library verilog;
use verilog.vl_types.all;
entity regfile_filter_sv_unit is
end regfile_filter_sv_unit;
