library verilog;
use verilog.vl_types.all;
entity control_sv_unit is
end control_sv_unit;
