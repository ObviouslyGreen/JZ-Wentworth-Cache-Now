library verilog;
use verilog.vl_types.all;
entity control_rom_sv_unit is
end control_rom_sv_unit;
