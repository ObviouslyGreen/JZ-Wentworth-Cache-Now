library verilog;
use verilog.vl_types.all;
entity mp2_sv_unit is
end mp2_sv_unit;
