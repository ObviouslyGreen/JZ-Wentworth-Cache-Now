library verilog;
use verilog.vl_types.all;
entity sext_sv_unit is
end sext_sv_unit;
