/*
 * Hazard detection unit
 */
import lc3b_types::*;

module hazard_detector
(
    input clk,
    input mem_read,
    input lc3b_opcode opcode,
    output logic bubble_enable
);

endmodule : hazard_detector
