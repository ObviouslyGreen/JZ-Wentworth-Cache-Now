library verilog;
use verilog.vl_types.all;
entity array_sv_unit is
end array_sv_unit;
