library verilog;
use verilog.vl_types.all;
entity ir_sv_unit is
end ir_sv_unit;
