library verilog;
use verilog.vl_types.all;
entity zext_sv_unit is
end zext_sv_unit;
