library verilog;
use verilog.vl_types.all;
entity zadj_sv_unit is
end zadj_sv_unit;
