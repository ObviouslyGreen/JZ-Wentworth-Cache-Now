library verilog;
use verilog.vl_types.all;
entity regfile_sv_unit is
end regfile_sv_unit;
