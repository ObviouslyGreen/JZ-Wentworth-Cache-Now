library verilog;
use verilog.vl_types.all;
entity stb_filter_sv_unit is
end stb_filter_sv_unit;
