library verilog;
use verilog.vl_types.all;
entity mp2_tb is
end mp2_tb;
