library verilog;
use verilog.vl_types.all;
entity adj_sv_unit is
end adj_sv_unit;
