library verilog;
use verilog.vl_types.all;
entity ctrl_register_sv_unit is
end ctrl_register_sv_unit;
