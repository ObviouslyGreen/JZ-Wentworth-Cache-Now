library verilog;
use verilog.vl_types.all;
entity datapath_sv_unit is
end datapath_sv_unit;
