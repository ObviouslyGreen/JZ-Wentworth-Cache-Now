library verilog;
use verilog.vl_types.all;
entity alu_sv_unit is
end alu_sv_unit;
