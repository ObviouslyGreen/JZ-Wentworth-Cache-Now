library verilog;
use verilog.vl_types.all;
entity mp3_tb is
end mp3_tb;
