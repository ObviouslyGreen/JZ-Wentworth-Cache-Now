library verilog;
use verilog.vl_types.all;
entity gencc_sv_unit is
end gencc_sv_unit;
