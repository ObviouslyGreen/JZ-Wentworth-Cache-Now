library verilog;
use verilog.vl_types.all;
entity byte_select_mux2_sv_unit is
end byte_select_mux2_sv_unit;
