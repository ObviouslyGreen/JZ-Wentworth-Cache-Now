library verilog;
use verilog.vl_types.all;
entity lc3b_types is
end lc3b_types;
