library verilog;
use verilog.vl_types.all;
entity data_membyte_filter_sv_unit is
end data_membyte_filter_sv_unit;
